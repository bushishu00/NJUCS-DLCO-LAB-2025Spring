`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/10/02 11:14:03
// Design Name: 
// Module Name: mul_32b
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mul_32b(
    output [63:0] p,         //�˻�
    output out_valid,        //�ߵ�ƽ��Чʱ����ʾ�˷�����������
    input clk,              //ʱ�� 
    input rst_n,             //��λ�źţ�����Ч
    input [31:0] x,           //������
    input [31:0] y,           //����
    input in_valid           //�ߵ�ƽ��Ч����ʾ�˷�����ʼ����
); 
//add your code here
endmodule
